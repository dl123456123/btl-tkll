module running_LED_v2(mode, mode_hz, auto, clk, reset, out, led7, led6, led5, led4, led3, led2, led1, led0, out_auto);
   input mode;
	input [2:0] mode_hz;
	input clk, reset, auto;
	output reg [25:0] out;
	output [6:0] led7, led6, led5, led4, led3, led2, led1, led0;
	output out_auto;
	reg temp;
	reg [3:0] auto_next=4'd0, count=4'd0;
	reg [3:0] mode_in=4'd0; 
	wire hz_led;
	wire hz_out;
	reg [2:0] countled=3'd0;
	reg [3:0] onled3210;
	wire [9:0] controlled54, controlled76;
	
	
	clock_divider c_d1(clk, mode_hz, hz_out);
	
	always @(posedge mode) begin
	   if(count<=4'd4) begin
		   count<=count+4'd1;
			if(count==4'd4) count<=4'd0;
		end
	end
	
	always @(*) begin
	   if(auto==1'b1) mode_in<=auto_next;
		else mode_in <= count;
	end
	
	always @(posedge hz_out, posedge reset) begin
	   if (reset) begin
		   out<=26'd0;
		end
		else begin
		   case(mode_in)
			4'd0: begin
			   case(out)
				26'b00000000000000000000000000: out<=26'b00000000000000000000000001;
				26'b00000000000000000000000001: out<=26'b00000000000000000000000010;
				26'b00000000000000000000000010: out<=26'b00000000000000000000000100;
				26'b00000000000000000000000100: out<=26'b00000000000000000000001000;
				26'b00000000000000000000001000: out<=26'b00000000000000000000010000;
				26'b00000000000000000000010000: out<=26'b00000000000000000000100000;
				26'b00000000000000000000100000: out<=26'b00000000000000000001000000;
				26'b00000000000000000001000000: out<=26'b00000000000000000010000000;
				26'b00000000000000000010000000: out<=26'b00000000000000000100000000;
				26'b00000000000000000100000000: out<=26'b00000000000000001000000000;
				26'b00000000000000001000000000: out<=26'b00000000000000010000000000;
				26'b00000000000000010000000000: out<=26'b00000000000000100000000000;
				26'b00000000000000100000000000: out<=26'b00000000000001000000000000;
				26'b00000000000001000000000000: out<=26'b00000000000010000000000000;
				26'b00000000000010000000000000: out<=26'b00000000000100000000000000;
				26'b00000000000100000000000000: out<=26'b00000000001000000000000000;
				26'b00000000001000000000000000: out<=26'b00000000010000000000000000;
				26'b00000000010000000000000000: out<=26'b00000000100000000000000000;
				26'b00000000100000000000000000: out<=26'b00000001000000000000000000;
				26'b00000001000000000000000000: out<=26'b00000010000000000000000000;
				26'b00000010000000000000000000: out<=26'b00000100000000000000000000;
				26'b00000100000000000000000000: out<=26'b00001000000000000000000000;
				26'b00001000000000000000000000: out<=26'b00010000000000000000000000;
				26'b00010000000000000000000000: out<=26'b00100000000000000000000000;
				26'b00100000000000000000000000: out<=26'b01000000000000000000000000;
				26'b01000000000000000000000000: out<=26'b10000000000000000000000000;
				26'b10000000000000000000000000: out<=26'b10000000000000000000000001;
				26'b10000000000000000000000001: out<=26'b10000000000000000000000010;
				26'b10000000000000000000000010: out<=26'b10000000000000000000000100;
				26'b10000000000000000000000100: out<=26'b10000000000000000000001000;
				26'b10000000000000000000001000: out<=26'b10000000000000000000010000;
				26'b10000000000000000000010000: out<=26'b10000000000000000000100000;
				26'b10000000000000000000100000: out<=26'b10000000000000000001000000;
				26'b10000000000000000001000000: out<=26'b10000000000000000010000000;
				26'b10000000000000000010000000: out<=26'b10000000000000000100000000;
				26'b10000000000000000100000000: out<=26'b10000000000000001000000000;
				26'b10000000000000001000000000: out<=26'b10000000000000010000000000;
				26'b10000000000000010000000000: out<=26'b10000000000000100000000000;
				26'b10000000000000100000000000: out<=26'b10000000000001000000000000;
				26'b10000000000001000000000000: out<=26'b10000000000010000000000000;
				26'b10000000000010000000000000: out<=26'b10000000000100000000000000;
				26'b10000000000100000000000000: out<=26'b10000000001000000000000000;
				26'b10000000001000000000000000: out<=26'b10000000010000000000000000;
				26'b10000000010000000000000000: out<=26'b10000000100000000000000000;
				26'b10000000100000000000000000: out<=26'b10000001000000000000000000;
				26'b10000001000000000000000000: out<=26'b10000010000000000000000000;
				26'b10000010000000000000000000: out<=26'b10000100000000000000000000;
				26'b10000100000000000000000000: out<=26'b10001000000000000000000000;
				26'b10001000000000000000000000: out<=26'b10010000000000000000000000;
				26'b10010000000000000000000000: out<=26'b10100000000000000000000000;
				26'b10100000000000000000000000: out<=26'b11000000000000000000000000;
				26'b11000000000000000000000000: out<=26'b11000000000000000000000001;
				26'b11000000000000000000000001: out<=26'b11000000000000000000000010;
				26'b11000000000000000000000010: out<=26'b11000000000000000000000100;
				26'b11000000000000000000000100: out<=26'b11000000000000000000001000;
				26'b11000000000000000000001000: out<=26'b11000000000000000000010000;
				26'b11000000000000000000010000: out<=26'b11000000000000000000100000;
				26'b11000000000000000000100000: out<=26'b11000000000000000001000000;
				26'b11000000000000000001000000: out<=26'b11000000000000000010000000;
				26'b11000000000000000010000000: out<=26'b11000000000000000100000000;
				26'b11000000000000000100000000: out<=26'b11000000000000001000000000;
				26'b11000000000000001000000000: out<=26'b11000000000000010000000000;
				26'b11000000000000010000000000: out<=26'b11000000000000100000000000;
				26'b11000000000000100000000000: out<=26'b11000000000001000000000000;
				26'b11000000000001000000000000: out<=26'b11000000000010000000000000;
				26'b11000000000010000000000000: out<=26'b11000000000100000000000000;
				26'b11000000000100000000000000: out<=26'b11000000001000000000000000;
				26'b11000000001000000000000000: out<=26'b11000000010000000000000000;
				26'b11000000010000000000000000: out<=26'b11000000100000000000000000;
				26'b11000000100000000000000000: out<=26'b11000001000000000000000000;
				26'b11000001000000000000000000: out<=26'b11000010000000000000000000;
				26'b11000010000000000000000000: out<=26'b11000100000000000000000000;
				26'b11000100000000000000000000: out<=26'b11001000000000000000000000;
				26'b11001000000000000000000000: out<=26'b11010000000000000000000000;
				26'b11010000000000000000000000: out<=26'b11100000000000000000000000;
				26'b11100000000000000000000000: out<=26'b11100000000000000000000001;
				26'b11100000000000000000000001: out<=26'b11100000000000000000000010;
				26'b11100000000000000000000010: out<=26'b11100000000000000000000100;
				26'b11100000000000000000000100: out<=26'b11100000000000000000001000;
				26'b11100000000000000000001000: out<=26'b11100000000000000000010000;
				26'b11100000000000000000010000: out<=26'b11100000000000000000100000;
				26'b11100000000000000000100000: out<=26'b11100000000000000001000000;
				26'b11100000000000000001000000: out<=26'b11100000000000000010000000;
				26'b11100000000000000010000000: out<=26'b11100000000000000100000000;
				26'b11100000000000000100000000: out<=26'b11100000000000001000000000;
				26'b11100000000000001000000000: out<=26'b11100000000000010000000000;
				26'b11100000000000010000000000: out<=26'b11100000000000100000000000;
				26'b11100000000000100000000000: out<=26'b11100000000001000000000000;
				26'b11100000000001000000000000: out<=26'b11100000000010000000000000;
				26'b11100000000010000000000000: out<=26'b11100000000100000000000000;
				26'b11100000000100000000000000: out<=26'b11100000001000000000000000;
				26'b11100000001000000000000000: out<=26'b11100000010000000000000000;
				26'b11100000010000000000000000: out<=26'b11100000100000000000000000;
				26'b11100000100000000000000000: out<=26'b11100001000000000000000000;
				26'b11100001000000000000000000: out<=26'b11100010000000000000000000;
				26'b11100010000000000000000000: out<=26'b11100100000000000000000000;
				26'b11100100000000000000000000: out<=26'b11101000000000000000000000;
				26'b11101000000000000000000000: out<=26'b11110000000000000000000000;
				26'b11110000000000000000000000: out<=26'b11110000000000000000000001;
				26'b11110000000000000000000001: out<=26'b11110000000000000000000010;
				26'b11110000000000000000000010: out<=26'b11110000000000000000000100;
				26'b11110000000000000000000100: out<=26'b11110000000000000000001000;
				26'b11110000000000000000001000: out<=26'b11110000000000000000010000;
				26'b11110000000000000000010000: out<=26'b11110000000000000000100000;
				26'b11110000000000000000100000: out<=26'b11110000000000000001000000;
				26'b11110000000000000001000000: out<=26'b11110000000000000010000000;
				26'b11110000000000000010000000: out<=26'b11110000000000000100000000;
				26'b11110000000000000100000000: out<=26'b11110000000000001000000000;
				26'b11110000000000001000000000: out<=26'b11110000000000010000000000;
				26'b11110000000000010000000000: out<=26'b11110000000000100000000000;
				26'b11110000000000100000000000: out<=26'b11110000000001000000000000;
				26'b11110000000001000000000000: out<=26'b11110000000010000000000000;
				26'b11110000000010000000000000: out<=26'b11110000000100000000000000;
				26'b11110000000100000000000000: out<=26'b11110000001000000000000000;
				26'b11110000001000000000000000: out<=26'b11110000010000000000000000;
				26'b11110000010000000000000000: out<=26'b11110000100000000000000000;
				26'b11110000100000000000000000: out<=26'b11110001000000000000000000;
				26'b11110001000000000000000000: out<=26'b11110010000000000000000000;
				26'b11110010000000000000000000: out<=26'b11110100000000000000000000;
				26'b11110100000000000000000000: out<=26'b11111000000000000000000000;
				26'b11111000000000000000000000: out<=26'b11111000000000000000000001;
				26'b11111000000000000000000001: out<=26'b11111000000000000000000010;
				26'b11111000000000000000000010: out<=26'b11111000000000000000000100;
				26'b11111000000000000000000100: out<=26'b11111000000000000000001000;
				26'b11111000000000000000001000: out<=26'b11111000000000000000010000;
				26'b11111000000000000000010000: out<=26'b11111000000000000000100000;
				26'b11111000000000000000100000: out<=26'b11111000000000000001000000;
				26'b11111000000000000001000000: out<=26'b11111000000000000010000000;
				26'b11111000000000000010000000: out<=26'b11111000000000000100000000;
				26'b11111000000000000100000000: out<=26'b11111000000000001000000000;
				26'b11111000000000001000000000: out<=26'b11111000000000010000000000;
				26'b11111000000000010000000000: out<=26'b11111000000000100000000000;
				26'b11111000000000100000000000: out<=26'b11111000000001000000000000;
				26'b11111000000001000000000000: out<=26'b11111000000010000000000000;
				26'b11111000000010000000000000: out<=26'b11111000000100000000000000;
				26'b11111000000100000000000000: out<=26'b11111000001000000000000000;
				26'b11111000001000000000000000: out<=26'b11111000010000000000000000;
				26'b11111000010000000000000000: out<=26'b11111000100000000000000000;
				26'b11111000100000000000000000: out<=26'b11111001000000000000000000;
				26'b11111001000000000000000000: out<=26'b11111010000000000000000000;
				26'b11111010000000000000000000: out<=26'b11111100000000000000000000;
				26'b11111100000000000000000000: out<=26'b11111100000000000000000001;
				26'b11111100000000000000000001: out<=26'b11111100000000000000000010;
				26'b11111100000000000000000010: out<=26'b11111100000000000000000100;
				26'b11111100000000000000000100: out<=26'b11111100000000000000001000;
				26'b11111100000000000000001000: out<=26'b11111100000000000000010000;
				26'b11111100000000000000010000: out<=26'b11111100000000000000100000;
				26'b11111100000000000000100000: out<=26'b11111100000000000001000000;
				26'b11111100000000000001000000: out<=26'b11111100000000000010000000;
				26'b11111100000000000010000000: out<=26'b11111100000000000100000000;
				26'b11111100000000000100000000: out<=26'b11111100000000001000000000;
				26'b11111100000000001000000000: out<=26'b11111100000000010000000000;
				26'b11111100000000010000000000: out<=26'b11111100000000100000000000;
				26'b11111100000000100000000000: out<=26'b11111100000001000000000000;
				26'b11111100000001000000000000: out<=26'b11111100000010000000000000;
				26'b11111100000010000000000000: out<=26'b11111100000100000000000000;
				26'b11111100000100000000000000: out<=26'b11111100001000000000000000;
				26'b11111100001000000000000000: out<=26'b11111100010000000000000000;
				26'b11111100010000000000000000: out<=26'b11111100100000000000000000;
				26'b11111100100000000000000000: out<=26'b11111101000000000000000000;
				26'b11111101000000000000000000: out<=26'b11111110000000000000000000;
				26'b11111110000000000000000000: out<=26'b11111110000000000000000001;
				26'b11111110000000000000000001: out<=26'b11111110000000000000000010;
				26'b11111110000000000000000010: out<=26'b11111110000000000000000100;
				26'b11111110000000000000000100: out<=26'b11111110000000000000001000;
				26'b11111110000000000000001000: out<=26'b11111110000000000000010000;
				26'b11111110000000000000010000: out<=26'b11111110000000000000100000;
				26'b11111110000000000000100000: out<=26'b11111110000000000001000000;
				26'b11111110000000000001000000: out<=26'b11111110000000000010000000;
				26'b11111110000000000010000000: out<=26'b11111110000000000100000000;
				26'b11111110000000000100000000: out<=26'b11111110000000001000000000;
				26'b11111110000000001000000000: out<=26'b11111110000000010000000000;
				26'b11111110000000010000000000: out<=26'b11111110000000100000000000;
				26'b11111110000000100000000000: out<=26'b11111110000001000000000000;
				26'b11111110000001000000000000: out<=26'b11111110000010000000000000;
				26'b11111110000010000000000000: out<=26'b11111110000100000000000000;
				26'b11111110000100000000000000: out<=26'b11111110001000000000000000;
				26'b11111110001000000000000000: out<=26'b11111110010000000000000000;
				26'b11111110010000000000000000: out<=26'b11111110100000000000000000;
				26'b11111110100000000000000000: out<=26'b11111111000000000000000000;
				26'b11111111000000000000000000: out<=26'b11111111000000000000000001;
				26'b11111111000000000000000001: out<=26'b11111111000000000000000010;
				26'b11111111000000000000000010: out<=26'b11111111000000000000000100;
				26'b11111111000000000000000100: out<=26'b11111111000000000000001000;
				26'b11111111000000000000001000: out<=26'b11111111000000000000010000;
				26'b11111111000000000000010000: out<=26'b11111111000000000000100000;
				26'b11111111000000000000100000: out<=26'b11111111000000000001000000;
				26'b11111111000000000001000000: out<=26'b11111111000000000010000000;
				26'b11111111000000000010000000: out<=26'b11111111000000000100000000;
				26'b11111111000000000100000000: out<=26'b11111111000000001000000000;
				26'b11111111000000001000000000: out<=26'b11111111000000010000000000;
				26'b11111111000000010000000000: out<=26'b11111111000000100000000000;
				26'b11111111000000100000000000: out<=26'b11111111000001000000000000;
				26'b11111111000001000000000000: out<=26'b11111111000010000000000000;
				26'b11111111000010000000000000: out<=26'b11111111000100000000000000;
				26'b11111111000100000000000000: out<=26'b11111111001000000000000000;
				26'b11111111001000000000000000: out<=26'b11111111010000000000000000;
				26'b11111111010000000000000000: out<=26'b11111111100000000000000000;
				26'b11111111100000000000000000: out<=26'b11111111100000000000000001;
				26'b11111111100000000000000001: out<=26'b11111111100000000000000010;
				26'b11111111100000000000000010: out<=26'b11111111100000000000000100;
				26'b11111111100000000000000100: out<=26'b11111111100000000000001000;
				26'b11111111100000000000001000: out<=26'b11111111100000000000010000;
				26'b11111111100000000000010000: out<=26'b11111111100000000000100000;
				26'b11111111100000000000100000: out<=26'b11111111100000000001000000;
				26'b11111111100000000001000000: out<=26'b11111111100000000010000000;
				26'b11111111100000000010000000: out<=26'b11111111100000000100000000;
				26'b11111111100000000100000000: out<=26'b11111111100000001000000000;
				26'b11111111100000001000000000: out<=26'b11111111100000010000000000;
				26'b11111111100000010000000000: out<=26'b11111111100000100000000000;
				26'b11111111100000100000000000: out<=26'b11111111100001000000000000;
				26'b11111111100001000000000000: out<=26'b11111111100010000000000000;
				26'b11111111100010000000000000: out<=26'b11111111100100000000000000;
				26'b11111111100100000000000000: out<=26'b11111111101000000000000000;
				26'b11111111101000000000000000: out<=26'b11111111110000000000000000;
				26'b11111111110000000000000000: out<=26'b11111111110000000000000001;
				26'b11111111110000000000000001: out<=26'b11111111110000000000000010;
				26'b11111111110000000000000010: out<=26'b11111111110000000000000100;
				26'b11111111110000000000000100: out<=26'b11111111110000000000001000;
				26'b11111111110000000000001000: out<=26'b11111111110000000000010000;
				26'b11111111110000000000010000: out<=26'b11111111110000000000100000;
				26'b11111111110000000000100000: out<=26'b11111111110000000001000000;
				26'b11111111110000000001000000: out<=26'b11111111110000000010000000;
				26'b11111111110000000010000000: out<=26'b11111111110000000100000000;
				26'b11111111110000000100000000: out<=26'b11111111110000001000000000;
				26'b11111111110000001000000000: out<=26'b11111111110000010000000000;
				26'b11111111110000010000000000: out<=26'b11111111110000100000000000;
				26'b11111111110000100000000000: out<=26'b11111111110001000000000000;
				26'b11111111110001000000000000: out<=26'b11111111110010000000000000;
				26'b11111111110010000000000000: out<=26'b11111111110100000000000000;
				26'b11111111110100000000000000: out<=26'b11111111111000000000000000;
				26'b11111111111000000000000000: out<=26'b11111111111000000000000001;
				26'b11111111111000000000000001: out<=26'b11111111111000000000000010;
				26'b11111111111000000000000010: out<=26'b11111111111000000000000100;
				26'b11111111111000000000000100: out<=26'b11111111111000000000001000;
				26'b11111111111000000000001000: out<=26'b11111111111000000000010000;
				26'b11111111111000000000010000: out<=26'b11111111111000000000100000;
				26'b11111111111000000000100000: out<=26'b11111111111000000001000000;
				26'b11111111111000000001000000: out<=26'b11111111111000000010000000;
				26'b11111111111000000010000000: out<=26'b11111111111000000100000000;
				26'b11111111111000000100000000: out<=26'b11111111111000001000000000;
				26'b11111111111000001000000000: out<=26'b11111111111000010000000000;
				26'b11111111111000010000000000: out<=26'b11111111111000100000000000;
				26'b11111111111000100000000000: out<=26'b11111111111001000000000000;
				26'b11111111111001000000000000: out<=26'b11111111111010000000000000;
				26'b11111111111010000000000000: out<=26'b11111111111100000000000000;
				26'b11111111111100000000000000: out<=26'b11111111111100000000000001;
				26'b11111111111100000000000001: out<=26'b11111111111100000000000010;
				26'b11111111111100000000000010: out<=26'b11111111111100000000000100;
				26'b11111111111100000000000100: out<=26'b11111111111100000000001000;
				26'b11111111111100000000001000: out<=26'b11111111111100000000010000;
				26'b11111111111100000000010000: out<=26'b11111111111100000000100000;
				26'b11111111111100000000100000: out<=26'b11111111111100000001000000;
				26'b11111111111100000001000000: out<=26'b11111111111100000010000000;
				26'b11111111111100000010000000: out<=26'b11111111111100000100000000;
				26'b11111111111100000100000000: out<=26'b11111111111100001000000000;
				26'b11111111111100001000000000: out<=26'b11111111111100010000000000;
				26'b11111111111100010000000000: out<=26'b11111111111100100000000000;
				26'b11111111111100100000000000: out<=26'b11111111111101000000000000;
				26'b11111111111101000000000000: out<=26'b11111111111110000000000000;
				26'b11111111111110000000000000: out<=26'b11111111111110000000000001;
				26'b11111111111110000000000001: out<=26'b11111111111110000000000010;
				26'b11111111111110000000000010: out<=26'b11111111111110000000000100;
				26'b11111111111110000000000100: out<=26'b11111111111110000000001000;
				26'b11111111111110000000001000: out<=26'b11111111111110000000010000;
				26'b11111111111110000000010000: out<=26'b11111111111110000000100000;
				26'b11111111111110000000100000: out<=26'b11111111111110000001000000;
				26'b11111111111110000001000000: out<=26'b11111111111110000010000000;
				26'b11111111111110000010000000: out<=26'b11111111111110000100000000;
				26'b11111111111110000100000000: out<=26'b11111111111110001000000000;
				26'b11111111111110001000000000: out<=26'b11111111111110010000000000;
				26'b11111111111110010000000000: out<=26'b11111111111110100000000000;
				26'b11111111111110100000000000: out<=26'b11111111111111000000000000;
				26'b11111111111111000000000000: out<=26'b11111111111111000000000001;
				26'b11111111111111000000000001: out<=26'b11111111111111000000000010;
				26'b11111111111111000000000010: out<=26'b11111111111111000000000100;
				26'b11111111111111000000000100: out<=26'b11111111111111000000001000;
				26'b11111111111111000000001000: out<=26'b11111111111111000000010000;
				26'b11111111111111000000010000: out<=26'b11111111111111000000100000;
				26'b11111111111111000000100000: out<=26'b11111111111111000001000000;
				26'b11111111111111000001000000: out<=26'b11111111111111000010000000;
				26'b11111111111111000010000000: out<=26'b11111111111111000100000000;
				26'b11111111111111000100000000: out<=26'b11111111111111001000000000;
				26'b11111111111111001000000000: out<=26'b11111111111111010000000000;
				26'b11111111111111010000000000: out<=26'b11111111111111100000000000;
				26'b11111111111111100000000000: out<=26'b11111111111111100000000001;
				26'b11111111111111100000000001: out<=26'b11111111111111100000000010;
				26'b11111111111111100000000010: out<=26'b11111111111111100000000100;
				26'b11111111111111100000000100: out<=26'b11111111111111100000001000;
				26'b11111111111111100000001000: out<=26'b11111111111111100000010000;
				26'b11111111111111100000010000: out<=26'b11111111111111100000100000;
				26'b11111111111111100000100000: out<=26'b11111111111111100001000000;
				26'b11111111111111100001000000: out<=26'b11111111111111100010000000;
				26'b11111111111111100010000000: out<=26'b11111111111111100100000000;
				26'b11111111111111100100000000: out<=26'b11111111111111101000000000;
				26'b11111111111111101000000000: out<=26'b11111111111111110000000000;
				26'b11111111111111110000000000: out<=26'b11111111111111110000000001;
				26'b11111111111111110000000001: out<=26'b11111111111111110000000010;
				26'b11111111111111110000000010: out<=26'b11111111111111110000000100;
				26'b11111111111111110000000100: out<=26'b11111111111111110000001000;
				26'b11111111111111110000001000: out<=26'b11111111111111110000010000;
				26'b11111111111111110000010000: out<=26'b11111111111111110000100000;
				26'b11111111111111110000100000: out<=26'b11111111111111110001000000;
				26'b11111111111111110001000000: out<=26'b11111111111111110010000000;
				26'b11111111111111110010000000: out<=26'b11111111111111110100000000;
				26'b11111111111111110100000000: out<=26'b11111111111111111000000000;
				26'b11111111111111111000000000: out<=26'b11111111111111111000000001;
				26'b11111111111111111000000001: out<=26'b11111111111111111000000010;
				26'b11111111111111111000000010: out<=26'b11111111111111111000000100;
				26'b11111111111111111000000100: out<=26'b11111111111111111000001000;
				26'b11111111111111111000001000: out<=26'b11111111111111111000010000;
				26'b11111111111111111000010000: out<=26'b11111111111111111000100000;
				26'b11111111111111111000100000: out<=26'b11111111111111111001000000;
				26'b11111111111111111001000000: out<=26'b11111111111111111010000000;
				26'b11111111111111111010000000: out<=26'b11111111111111111100000000;
				26'b11111111111111111100000000: out<=26'b11111111111111111100000001;
				26'b11111111111111111100000001: out<=26'b11111111111111111100000010;
				26'b11111111111111111100000010: out<=26'b11111111111111111100000100;
				26'b11111111111111111100000100: out<=26'b11111111111111111100001000;
				26'b11111111111111111100001000: out<=26'b11111111111111111100010000;
				26'b11111111111111111100010000: out<=26'b11111111111111111100100000;
				26'b11111111111111111100100000: out<=26'b11111111111111111101000000;
				26'b11111111111111111101000000: out<=26'b11111111111111111110000000;
				26'b11111111111111111110000000: out<=26'b11111111111111111110000001;
				26'b11111111111111111110000001: out<=26'b11111111111111111110000010;
				26'b11111111111111111110000010: out<=26'b11111111111111111110000100;
				26'b11111111111111111110000100: out<=26'b11111111111111111110001000;
				26'b11111111111111111110001000: out<=26'b11111111111111111110010000;
				26'b11111111111111111110010000: out<=26'b11111111111111111110100000;
				26'b11111111111111111110100000: out<=26'b11111111111111111111000000;
				26'b11111111111111111111000000: out<=26'b11111111111111111111000001;
				26'b11111111111111111111000001: out<=26'b11111111111111111111000010;
				26'b11111111111111111111000010: out<=26'b11111111111111111111000100;
				26'b11111111111111111111000100: out<=26'b11111111111111111111001000;
				26'b11111111111111111111001000: out<=26'b11111111111111111111010000;
				26'b11111111111111111111010000: out<=26'b11111111111111111111100000;
				26'b11111111111111111111100000: out<=26'b11111111111111111111100001;
				26'b11111111111111111111100001: out<=26'b11111111111111111111100010;
				26'b11111111111111111111100010: out<=26'b11111111111111111111100100;
				26'b11111111111111111111100100: out<=26'b11111111111111111111101000;
				26'b11111111111111111111101000: out<=26'b11111111111111111111110000;
				26'b11111111111111111111110000: out<=26'b11111111111111111111110001;
				26'b11111111111111111111110001: out<=26'b11111111111111111111110010;
				26'b11111111111111111111110010: out<=26'b11111111111111111111110100;
				26'b11111111111111111111110100: out<=26'b11111111111111111111111000;
				26'b11111111111111111111111000: out<=26'b11111111111111111111111001;
				26'b11111111111111111111111001: out<=26'b11111111111111111111111010;
				26'b11111111111111111111111010: out<=26'b11111111111111111111111100;
				26'b11111111111111111111111100: out<=26'b11111111111111111111111101;
				26'b11111111111111111111111101: out<=26'b11111111111111111111111110;
				26'b11111111111111111111111110: out<=26'b11111111111111111111111111;
				26'b11111111111111111111111111: begin
				   out<=26'b00000000000000000000000000;
					auto_next<=4'd1;
				end
				default: out<=26'b00000000000000000000000000;
				endcase
         end
			4'd1: begin
			   case({temp,out})
			   27'b000000000000000000000000000: {temp,out}<=27'b000000000000000000000000001;
				27'b000000000000000000000000001: {temp,out}<=27'b000000000000000000000000011;
				27'b000000000000000000000000011: {temp,out}<=27'b000000000000000000000000111;
				27'b000000000000000000000000111: {temp,out}<=27'b000000000000000000000001111;
				27'b000000000000000000000001111: {temp,out}<=27'b000000000000000000000011111;
				27'b000000000000000000000011111: {temp,out}<=27'b000000000000000000000101111;
				27'b000000000000000000000101111: {temp,out}<=27'b000000000000000000001010111;
				27'b000000000000000000001010111: {temp,out}<=27'b000000000000000000010101011;
				27'b000000000000000000010101011: {temp,out}<=27'b000000000000000000101010101;
				27'b000000000000000000101010101: {temp,out}<=27'b000000000000000001010101010;
				27'b000000000000000001010101010: {temp,out}<=27'b000000000000000010101010100;
				27'b000000000000000010101010100: {temp,out}<=27'b000000000000000101010101000;
				27'b000000000000000101010101000: {temp,out}<=27'b000000000000001010101010000;
				27'b000000000000001010101010000: {temp,out}<=27'b000000000000010101010100000;
				27'b000000000000010101010100000: {temp,out}<=27'b000000000000101010101000000;
				27'b000000000000101010101000000: {temp,out}<=27'b000000000001010101010000000;
				27'b000000000001010101010000000: {temp,out}<=27'b000000000010101010100000000;
				27'b000000000010101010100000000: {temp,out}<=27'b000000000101010101000000000;
				27'b000000000101010101000000000: {temp,out}<=27'b000000001010101010000000000;
				27'b000000001010101010000000000: {temp,out}<=27'b000000010101010100000000000;
				27'b000000010101010100000000000: {temp,out}<=27'b000000101010101000000000000;
				27'b000000101010101000000000000: {temp,out}<=27'b000001010101010000000000000;
				27'b000001010101010000000000000: {temp,out}<=27'b000010101010100000000000000;
				27'b000010101010100000000000000: {temp,out}<=27'b000101010101000000000000000;
				27'b000101010101000000000000000: {temp,out}<=27'b001010101010000000000000000;
				27'b001010101010000000000000000: {temp,out}<=27'b010101010100000000000000000;
				27'b010101010100000000000000000: {temp,out}<=27'b011010101000000000000000000;
				27'b011010101000000000000000000: {temp,out}<=27'b011101010000000000000000000;
				27'b011101010000000000000000000: {temp,out}<=27'b011110100000000000000000000;
				27'b011110100000000000000000000: {temp,out}<=27'b011111000000000000000000000;
				27'b011111000000000000000000000: {temp,out}<=27'b111110100000000000000000000;
				27'b111110100000000000000000000: {temp,out}<=27'b111101010000000000000000000;
				27'b111101010000000000000000000: {temp,out}<=27'b111010101000000000000000000;
				27'b111010101000000000000000000: {temp,out}<=27'b110101010100000000000000000;
				27'b110101010100000000000000000: {temp,out}<=27'b101010101010000000000000000;
				27'b101010101010000000000000000: {temp,out}<=27'b100101010101000000000000000;
				27'b100101010101000000000000000: {temp,out}<=27'b100010101010100000000000000;
				27'b100010101010100000000000000: {temp,out}<=27'b100001010101010000000000000;
				27'b100001010101010000000000000: {temp,out}<=27'b100000101010101000000000000;
				27'b100000101010101000000000000: {temp,out}<=27'b100000010101010100000000000;
				27'b100000010101010100000000000: {temp,out}<=27'b100000001010101010000000000;
				27'b100000001010101010000000000: {temp,out}<=27'b100000000101010101000000000;
				27'b100000000101010101000000000: {temp,out}<=27'b100000000010101010100000000;
				27'b100000000010101010100000000: {temp,out}<=27'b100000000001010101010000000;
				27'b100000000001010101010000000: {temp,out}<=27'b100000000000101010101000000;
				27'b100000000000101010101000000: {temp,out}<=27'b100000000000010101010100000;
				27'b100000000000010101010100000: {temp,out}<=27'b100000000000001010101010000;
				27'b100000000000001010101010000: {temp,out}<=27'b100000000000000101010101000;
				27'b100000000000000101010101000: {temp,out}<=27'b100000000000000010101010100;
				27'b100000000000000010101010100: {temp,out}<=27'b100000000000000001010101010;
				27'b100000000000000001010101010: {temp,out}<=27'b100000000000000000101010101;
				27'b100000000000000000101010101: {temp,out}<=27'b100000000000000000010101011;
				27'b100000000000000000010101011: {temp,out}<=27'b100000000000000000001010111;
				27'b100000000000000000001010111: {temp,out}<=27'b100000000000000000000101111;
				27'b100000000000000000000101111: begin
				   {temp,out}<=27'b100000000000000000000011111;
					auto_next<=4'd2;
				end
				27'b100000000000000000000011111: {temp,out}<=27'b000000000000000000000101111;
				default: {temp,out}<=27'b00000000000000000000000000;
				endcase
			end
			4'd2: begin
			   case({temp,out})
				27'b000000000000000000000000000: {temp,out}<=27'b000000000000000000000000001;
				27'b000000000000000000000000001: {temp,out}<=27'b000000000000000000000000010;
				27'b000000000000000000000000010: {temp,out}<=27'b000000000000000000000000100;
				27'b000000000000000000000000100: {temp,out}<=27'b000000000000000000000001000;
				27'b000000000000000000000001000: {temp,out}<=27'b000000000000000000000010000;
				27'b000000000000000000000010000: {temp,out}<=27'b000000000000000000000100000;
				27'b000000000000000000000100000: {temp,out}<=27'b000000000000000000001000000;
				27'b000000000000000000001000000: {temp,out}<=27'b000000000000000000010000000;
				27'b000000000000000000010000000: {temp,out}<=27'b000000000000000000100000000;
				27'b000000000000000000100000000: {temp,out}<=27'b000000000000000001000000000;
				27'b000000000000000001000000000: {temp,out}<=27'b000000000000000010000000000;
				27'b000000000000000010000000000: {temp,out}<=27'b000000000000000100000000000;
				27'b000000000000000100000000000: {temp,out}<=27'b000000000000001000000000000;
				27'b000000000000001000000000000: {temp,out}<=27'b000000000000111100000000000;
			   27'b000000000000111100000000000: {temp,out}<=27'b100000000000111100000000000;
				27'b100000000000111100000000000: {temp,out}<=27'b000000000010111101000000000;
				27'b000000000010111101000000000: {temp,out}<=27'b100000000010111101000000000;
				27'b100000000010111101000000000: {temp,out}<=27'b000000001010111101010000000;
				27'b000000001010111101010000000: {temp,out}<=27'b100000001010111101010000000;
				27'b100000001010111101010000000: {temp,out}<=27'b000000101010111101010100000;
				27'b000000101010111101010100000: {temp,out}<=27'b100000101010111101010100000;
				27'b100000101010111101010100000: {temp,out}<=27'b000010101010111101010101000;
				27'b000010101010111101010101000: {temp,out}<=27'b100010101010111101010101000;
				27'b100010101010111101010101000: {temp,out}<=27'b001010101010111101010101010;
				27'b001010101010111101010101010: {temp,out}<=27'b101010101010111101010101010;
				27'b101010101010111101010101010: {temp,out}<=27'b001010101010100101010101010;
				27'b001010101010100101010101010: {temp,out}<=27'b001010101010000001010101010;
				27'b001010101010000001010101010: {temp,out}<=27'b001010101000000000010101010;
				27'b001010101000000000010101010: {temp,out}<=27'b001010100000000000000101010;
				27'b001010100000000000000101010: {temp,out}<=27'b001010000000000000000001010;
				27'b001010000000000000000001010: {temp,out}<=27'b001000000000000000000000010;
				27'b001000000000000000000000010: begin
				   {temp,out}<=27'b000000000000000000000000000;
					auto_next<=4'd3;
				end
				default: {temp,out}<=27'b000000000000000000000000000;
				endcase
			end
			4'd3: begin
			   case(out)
				26'b00000000000000000000000000: out<=26'b00000000000000000000000001;
				26'b00000000000000000000000001: out<=26'b00000000000000000000110001;
				26'b00000000000000000000110001: out<=26'b00010000000000000000110001;
				26'b00010000000000000000110001: out<=26'b00010000000111000000110001;
				26'b00010000000111000000110001: out<=26'b00010011000111000000110001;
				26'b00010011000111000000110001: out<=26'b00010011000111001100110001;
				26'b00010011000111001100110001: out<=26'b11010011000111001100110001;
				26'b11010011000111001100110001: out<=26'b11010011000111001100111111;
				26'b11010011000111001100111111: out<=26'b11010011101111001100111111;
            26'b11010011101111001100111111: out<=26'b11010011101111001110111111;
            26'b11010011101111001110111111: out<=26'b11011011101111001110111111;
            26'b11011011101111001110111111: out<=26'b11011011101111101110111111;
            26'b11011011101111101110111111: out<=26'b11111011101111101110111111;
            26'b11111011101111101110111111: out<=26'b11111011111111101110111111;
	         26'b11111011111111101110111111: out<=26'b11111011111111111110111111;
		      26'b11111011111111111110111111: out<=26'b11111011111111111111111111;
			   26'b11111011111111111111111111: out<=26'b11111111111111111111111111;
				26'b11111111111111111111111111: begin
				   out<=26'b00000000000000000000000000;
					auto_next<=4'd0;
				end
				default: out<=26'b00000000000000000000000000;
				endcase
			end
		   default: out<=26'b11111111111111111111111111;
			endcase
		end
	end
	
	clock_divider c_d2(clk, 3'd2, hz_led);
	
	always @(posedge hz_led) begin
	   if(countled<=3'd5) begin
		   countled<=countled+3'd1;
			if(countled>=3'd0 && countled<=3'd3) onled3210[countled]<=1'b1;
		end
		if(countled==3'd6) begin
		   countled<=3'd0;
			onled3210<=4'd0;
		end
	end
	
	led7_decoder l3(onled3210[0], 4'b1110, led3);
	led7_decoder l2(onled3210[1], 4'b1111, led2);
	led7_decoder l1(onled3210[2], 4'b0001, led1);
	led7_decoder l0(onled3210[3], 4'b1001, led0);
	
	assign controlled76[8:5]=mode_in/4'd10;
	assign controlled76[3:0]=mode_in%4'd10;
	assign controlled76[9]=(controlled76[8:5]==4'd0)? 1'b0:1'b1;
	assign controlled76[4]=1'b1;
	
	led7_decoder l7(controlled76[9], controlled76[8:5], led7);
	led7_decoder l6(controlled76[4], controlled76[3:0], led6);
	
	assign controlled54=(mode_hz==3'd0)? 10'b1000010101:
	                    (mode_hz==3'd1)? 10'b0000010001:
							  (mode_hz==3'd2)? 10'b0000010010:
							  (mode_hz==3'd3)? 10'b0000010100:
							  (mode_hz==3'd4)? 10'b0000011000:10'b0000011000;
							 
	led7_decoder l5(controlled54[9], controlled54[8:5], led5);
	led7_decoder l4(controlled54[4], controlled54[3:0], led4);
	
	assign out_auto=auto;
	
endmodule
	